module rom(addr,data);
input [3:0] addr;
output reg [11:0] data;

always@ (*)
    case(addr)
        
        4'b0001 : data = 12'b000001100000; // 1
        4'b0010 : data = 12'b111000100000; // 2
        4'b0011 : data = 12'b100000100000; // 3 
        4'b0100 : data = 12'b110000101100; // 4
        4'b0101 : data = 12'b110101000100; // 5
        4'b0110 : data = 12'b111101010000; // 6
        4'b0111 : data = 12'b000100001001; // 7
        4'b1000 : data = 12'b001000000001; // 8
        4'b1001 : data = 12'b001000000100; // 9
        4'b1010 : data = 12'b010001000100; // a
        4'b1011 : data = 12'b010101100000; // b
        4'b1100 : data = 12'b011111000100; // c
        4'b1101 : data = 12'b100100100000; // d
        4'b1110 : data = 12'b101010001000; // e
        default : data = 12'b101100100000; // f
    endcase 

endmodule