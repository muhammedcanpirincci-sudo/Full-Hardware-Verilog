
module decoder8bit(enRAM, address, out);
input enRAM;
input [7:0] address;
output reg [255:0] out ;

always@(enRAM or address)begin
out = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	if(enRAM == 1'b1)
		begin
			out[address] = 1'b1;
		end 
end
endmodule